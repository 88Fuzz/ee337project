// $Id: $
// File name:   AES.sv
// Created:     12/1/2013
// Author:      Josh Nichols
// Lab Section: 002
// Version:     1.0  Initial Design Entry
// Description: Top Level Wrapper

module AES
(
  input wire HCLK,
  input wire HNRST,
	input wire clk,
	input wire n_rst,
	input wire [31:0] HADDR,
	input wire [2:0] HBURST,
	input wire HMASTLOCK,
	input wire [3:0] HPORT,
	input wire [2:0] HSIZE,
	input wire [1:0] HTRANS,
	input wire [127:0] HWDATA,
	input wire HWRITE,
	input wire HSELx,
	input wire HREADY,
	input wire sramBigDumpNum,
	input wire sramBigDump,
	output reg HRESP,
	output reg [127:0] HRDATA,
	output reg HREADYOUT
);







//top level sram signals
wire sramBigReadEnable;
wire sramBigWriteEnable;
wire [127:0]sramBigWriteValue;
reg [127:0]sramBigReadValue;
wire [15:0]sramBigAddr;
//wire sramBigDump;//////////////////////////////////////////////////////////////
//wire [2:0]sramBigDumpNum;
wire [2:0]sramBigInitNum;
wire sramBigInit;

//assign sramBigDumpNum=0;////////////////
//assign sramBigInitNum=0;

//keyexpansion sram signals
wire [127:0]sramWriteValue_keyexp;
wire sramRead_keyexp;
wire sramWrite_keyexp;
wire sramDump_keyexp;
wire sramInit_keyexp;
wire [15:0]sramAddr_keyexp;
wire [2:0]sramDumpNum_keyexp;
wire [2:0]sramInitNum_keyexp;

assign sramDumpNum_keyexp=0;
assign sramInitNum_keyexp=0;


//aroundwrap sram signals		
wire sramWrite_around;
wire sramRead_around;
wire [15:0]sramAddr_around;
wire sramDump_around;
wire [2:0]sramDumpNum_around;
wire [2:0]sramInitNum_around;
wire sramInit_around;
wire [127:0]sramWriteValue_around;

assign sramDumpNum_around=0;
assign sramInitNum_around=0;

//sbyteswrap sram signals
wire sramWrite_sbytes;
wire sramRead_sbytes;
wire [15:0]sramAddr_sbytes;
wire sramDump_sbytes;
wire [2:0]sramDumpNum_sbytes;
wire [2:0]sramInitNum_sbytes;
wire sramInit_sbytes;
wire [127:0]sramWriteValue_sbytes;

assign sramDumpNum_sbytes=0;
assign sramInitNum_sbytes=0;

//mixcolumn sram signals
wire sramWrite_mcol;
wire sramRead_mcol;
wire [15:0]sramAddr_mcol;
wire sramDump_mcol;
wire [2:0]sramDumpNum_mcol;
wire [2:0]sramInitNum_mcol;
wire sramInit_mcol;
wire [127:0]sramWriteValue_mcol;

assign sramDumpNum_mcol=0;
assign sramInitNum_mcol=0;

//srows sram signals
wire sramWrite_srows;
wire sramRead_srows;
wire [15:0]sramAddr_srows;
wire sramDump_srows;
wire [2:0]sramDumpNum_srows;
wire [2:0]sramInitNum_srows;
wire sramInit_srows;
wire [127:0]sramWriteValue_srows;

assign sramDumpNum_srows=0;
assign sramInitNum_srows=0;


//wire [31:0]HADDR;
//wire [2:0]HBURST;
//wire HMASTLOCK;
//wire [3:0] HPORT;
//wire [2:0] HSIZE;
//wire [1:0] HTRANS;
//wire HWRITE;//high=write, low=read
//wire HSELx;
//wire HREADY;
wire addrMatch;
wire mWrite;
wire mRead;
wire dataReady;
wire invalid;



wire readk_enable;//master writing key
wire read_enable;//master writing data
wire write_enable;//master reading data
wire hready_enable;
//AMBA_inout sram signals
wire [127:0]sramWriteValue_AMBA;
wire sramRead_AMBA;
wire sramWrite_AMBA;
wire [15:0]sramAddr_AMBA;
wire sramDump_ADDR;
wire [2:0]sramDumpNum_AMBA;
wire [2:0]sramInitNum_AMBA;
wire sramInit_AMBA;



wire [3:0]roundnum;
wire hresp_error;
wire HCLK_fall;
wire HCLK_rise;




//assign sramBigDump=0;/////////////////////////////////////////////////////////////////////////////////////////////////////
//assign sramBigDumpNum=0;
assign sramBigInitNum=0;
assign sramBigInit=0;
assign sramBigAddr=sramAddr_AMBA|sramAddr_srows|sramAddr_mcol|sramAddr_sbytes|sramAddr_around|sramAddr_keyexp;
assign sramBigReadEnable=sramRead_AMBA|sramRead_srows|sramRead_mcol|sramRead_sbytes|sramRead_around|sramRead_keyexp;
assign sramBigWriteEnable=sramWrite_AMBA|sramWrite_srows|sramWrite_mcol|sramWrite_sbytes|sramWrite_around|sramWrite_keyexp;
assign sramBigWriteValue=sramWriteValue_AMBA|sramWriteValue_srows|sramWriteValue_mcol|sramWriteValue_sbytes|sramWriteValue_around|sramWriteValue_keyexp;


	controller controller
	(
		.clk(clk),
		.n_rst(n_rst),
		.addrMatch(addrMatch),
		.HSELx(HSELx),
		.mWrite(mWrite),
		.dataReady(dataReady),
		.mRead(mRead),
		.keyexp_finished(keyexp_finished),
		.sbytes_finished(sbytes_finished),
		.srows_finished(srows_finished),
		.mcol_finished(mcol_finished),
		.around_finished(around_finished),
		.invalid(invalid),
		.HREADYOUT(hready_enable),
		.readk_enable(readk_enable),
		.read_enable(read_enable),
		.write_enable(write_enable),
		.keyexp_enable(keyexp_enable),
		.sbytes_enable(sbytes_enable),
		.srows_enable(srows_enable),
		.mcol_enable(mcol_enable),
		.around_enable(around_enable),
		.hresp_error(hresp_error),
		.roundnum(roundnum)
	);
	
	


	keyExpansion keyExpansion
	(
	  //INPUTS
		.clk(clk),
  		.n_rst(n_rst),
  		.roundNum(roundnum),
  		.enable(keyexp_enable),
  		.sramReadValue(sramBigReadValue),
  		//OUTPUTS
  		.expansionDone(keyexp_finished),
  		.sramWriteValue(sramWriteValue_keyexp),
  		.sramRead(sramRead_keyexp),
  		.sramWrite(sramWrite_keyexp),
  		.sramDump(sramDump_keyexp),
  		.sramInit(sramInit_keyexp),
  		.sramAddr(sramAddr_keyexp),
  		.sramDumpNum(sramDumpNum_keyexp),
  		.sramInitNum(sramInitNum_keyexp)
	);


  sbyteswrap sbyteswrap
  (
	.clk(clk),
  .n_rst(n_rst),
  .sbytes_enable(sbytes_enable),
  .sbytes_finished(sbytes_finished),
  .sramread_data(sramBigReadValue),
	.sramwrite_data(sramWriteValue_sbytes),
  .sramread(sramRead_sbytes),
  .sramwrite(sramWrite_sbytes),
  .sramdump(sramDump_sbytes),
  .sraminit(sramInit_sbytes),
  .sramaddr(sramAddr_sbytes),
  .sramdumpnum(sramDumpNum_sbytes),
  .sraminitnum(sramInitNum_sbytes)
  );	

/*	sbyteswrap sbyteswrap
	(
	  //INPUTES
		.clk(clk),
		.n_rst(n_rst),
		.sbytes_enable(sbytes_enable),
sramBigReadValue),
		//OUTPUTS
sramWrite_sbytes),
sramRead_sbytes),
sramAddr_sbytes),
sramDump_sbytes),
sramDumpNum_sbytes),
sramInitNum_sbytes),
sramInit_sbytes),
sramWriteValue_sbytes),
		.sbytes_finished(sbytes_finished)
	);*/




	mixcol mixcol
	(
	  //INPUT
	  .clk(clk),
	  .n_rst(n_rst),
		.mixcol_enable(mcol_enable),
    .sramReadValue(sramBigReadValue),
		//OUTPUT
    .sramWrite(sramWrite_mcol),
    .sramRead(sramRead_mcol),
    .sramAddr(sramAddr_mcol),
    .sramDump(sramDump_mcol),
    .sramDumpNum(sramDumpNum_mcol),
    .sramInitNum(sramInitNum_mcol),
    .sramInit(sramInit_mcol),
    .sramWriteValue(sramWriteValue_mcol),
		.mixcol_finished(mcol_finished)
	);
	
	


	srows srows
	(
	  //INPUT
	  .clk(clk),
	  .n_rst(n_rst),
	  .srows_enable(srows_enable),
    .sramReadValue(sramBigReadValue),
	  //OUTPUT
    .sramWrite(sramWrite_srows),
    .sramRead(sramRead_srows),
    .sramAddr(sramAddr_srows),
    .sramDump(sramDump_srows),
    .sramDumpNum(sramDumpNum_srows),
    .sramInitNum(sramInitNum_srows),
    .sramInit(sramInit_srows),
    .sramWriteValue(sramWriteValue_srows),
	  .srows_finished(srows_finished)
	);

	aroundwrap aroundwrap
	(
	  //INPUTS
		.clk(clk),
		.n_rst(n_rst),
		.around_enable(around_enable),
    .sramread_data(sramBigReadValue),		
		//OUTPUTS
    .sramwrite(sramWrite_around),
    .sramread(sramRead_around),
    .sramaddr(sramAddr_around),
    .sramdump(sramDump_around),
    .sramdumpnum(sramDumpNum_around),
    .sraminitnum(sramInitNum_around),
    .sraminit(sramInit_around),
    .sramwrite_data(sramWriteValue_around),
		.around_finished(around_finished)
	);
  
	AMBAsensor AMBAsensor
 (
  .HADDR(HADDR),
  .HBURST(HBURST),
  .HMASTLOCK(HMASTLOCK),
  .HPORT(HPORT),
  .HSIZE(HSIZE),
  .HTRANS(HTRANS),
  .HWRITE(HWRITE),//high=write, low=read
  .HSELx(HSELx),
  .HREADY(HREADY),
  .addrMatch(addrMatch),
  .mWrite(mWrite),
  .mRead(mRead),
  .dataReady(dataReady),
  .invalid(invalid)
 );
 
  HCLK_edgedet HCK_edgedet
(
  .clk(clk),
  .n_rst(n_rst),
  .HCLK(HCLK),
  .HCLK_rise(HCLK_rise),
  .HCLK_fall(HCLK_fall)
);


  AMBA_inout AMBA_inout
  (
  .HCLK(HCLK),
  .HNRST(HNRST),
  .HCLK_fall(HCLK_fall),
  .HCLK_rise(HCLK_rise),
  .clk(clk),
  .n_rst(n_rst),
  .writek_enable(readk_enable),//master writing key
  .writed_enable(read_enable),//master writing data
  .readd_enable(write_enable),//master reading data
  .hresp_error(hresp_error),
  .hready_enable(hready_enable),
  .read_data(sramBigReadValue),
  .HWDATA(HWDATA),
  .HRDATA(HRDATA),
  .write_data(sramWriteValue_AMBA),
  .HREADYOUT(HREADYOUT),
  .HRESP(HRESP),
  .read(sramRead_AMBA),
  .write(sramWrite_AMBA),
  .addr(sramAddr_AMBA),
  .dump(sramDump_ADDR),
  .dumpNum(sramDumpNum_AMBA),
  .initNum(sramInitNum_AMBA),
  .init(sramInit_AMBA)
  );


  testing_sram testing_sram
  (
  .read(sramBigReadEnable),
  .write(sramBigWriteEnable),
  .addr(sramBigAddr),
  .dump(sramBigDump),
  .dumpNum(sramBigDumpNum),
  .initNum(sramBigInitNum),
  .init(sramBigInit),
  .write_data(sramBigWriteValue),
  .read_data(sramBigReadValue)
  );
  
endmodule