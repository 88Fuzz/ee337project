library verilog;
use verilog.vl_types.all;
entity tb_flex_pts_sr is
end tb_flex_pts_sr;
