library verilog;
use verilog.vl_types.all;
entity tb_parallel_to_parallel is
end tb_parallel_to_parallel;
