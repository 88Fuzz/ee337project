module tb_flex_counter();

endmodule
