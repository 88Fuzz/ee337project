// $Id: $
// File name:   srows.sv
// Created:     11/18/2013
// Author:      Josh Nichols
// Lab Section: 002
// Version:     1.0  Initial Design Entry
// Description: Shift Rows

module srows
(
	input wire clk,
	input wire n_rst,
	input wire [127:0] sramReadValue,
	input wire srows_enable,
	output reg srows_finished,
	output reg [127:0] sramWriteValue,
	output reg sramRead,
	output reg sramWrite,
	output reg sramDump,
	output reg sramInit,
	output reg [15:0] sramAddr,
	output reg [2:0] sramDumpNum,
	output reg [2:0] sramInitNum
);
	reg [127:0] olddata;
	reg [127:0] newdata;
	reg [127:0] nextdata;
	reg [127:0] currdata;
	reg activate;
	reg currfinish;
	reg nextfinish;
	reg rstnextdata;

	typedef enum bit [3:0] {setaddr, idle, readsram1, readagain, shifter, writeaddr, writesram, finito, buff1, buff2} stateType;
	stateType state, nextstate;

	always@(posedge clk, negedge n_rst) begin
		if(n_rst == 1'b0) begin
			state <= idle;
			currfinish <= 0;
			currdata <= 0;
		end else begin
			state <= nextstate;
			currfinish <= nextfinish;
			currdata <= nextdata;
		end
	end

	assign olddata = sramReadValue;
	assign sramWriteValue = newdata;
	assign srows_finished = currfinish;

	always@(state, srows_enable) begin
		nextstate = state;
		case(state)
			idle: begin
				if(srows_enable) begin
					nextstate = setaddr;
				end else begin
					nextstate = idle;
				end
			end
			setaddr: begin
				nextstate = readsram1;
			end
			readsram1: begin
				nextstate = readagain;
			end
			readagain: begin
				nextstate = shifter;
			end
			shifter: begin
				nextstate = writeaddr;
			end
			writeaddr: begin
				nextstate = writesram;
			end
			writesram: begin
				nextstate = finito;
			end
			finito: begin
				nextstate = buff1;
			end
			buff1: begin
				nextstate = buff2;
			end
			buff2: begin
				nextstate = idle;
			end
			default: begin
				nextstate = state;
			end
		endcase
	end

	always@(state) begin
		//sramWriteValue = 1'b0;
		sramRead = 0;
		sramWrite = 0;
		sramDump = 0;
		sramInit = 0;
		sramAddr = 0;
		sramDumpNum = 0;
		sramInitNum = 0;
		nextfinish = 1'b0;
		activate = 1'b0;
		rstnextdata=0;
		case(state)
			idle: begin
			end
			setaddr: begin
				sramAddr = 32;
			end
			readsram1: begin
				sramAddr = 32;
				sramRead = 1'b1;
			end
			readagain: begin
			end
			shifter: begin
				activate = 1'b1;
			end
			writeaddr: begin
				sramAddr = 32;
			end
			writesram: begin
				sramAddr = 32;
				sramWrite = 1'b1;
			end
			finito: begin
				nextfinish = 1'b1;
				rstnextdata=1;
			end
			buff1: begin
			end
			buff2: begin
			end
			default: begin
			end
		endcase
	end

	assign newdata = currdata;

	//assign nextdata = activate ? {olddata[127:96],olddata[87:64],olddata[95:88],olddata[47:32],olddata[63:48],olddata[7:0],olddata[31:8]} : currdata;
	
	assign nextdata = rstnextdata ? 0 : activate ? {olddata[127:120],olddata[87:80],olddata[47:40],olddata[7:0],
	                              olddata[95:88],olddata[55:48],olddata[15:8],olddata[103:96],
	                              olddata[63:56],olddata[23:16],olddata[111:104],olddata[71:64],
	                              olddata[31:24],olddata[119:112],olddata[79:72],olddata[39:32]} : currdata;
	                              

//	assign srows_finished = (newdata == olddata) ? 1'b0 : 1'b1;
/*
	always@(posedge clk, negedge n_rst) begin
		if(n_rst == 1'b0) begin
			newdata <= olddata;
		end else begin
			if(srows_enable) begin
				newdata <= {olddata[31:0],olddata[63:40],olddata[39:32],olddata[95:80],olddata[79:64],olddata[127:119],olddata[119:96]};
				srows_finished = 1'b1;
			end
		end
	end		
*/

endmodule
