module HCLK_edgedet
(
);